pBAV       0� �� $  @  ����_��@�  ����������@�  ����������@�  ����������@�  ��������u��@�  ����������@�  ����������@�  ����������@�  ����������@�  ����������@�  ����������@�  ����������@�  ��������u��@�  ����������@�  ����������@�  ����������@�  ����������@�  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  �������� }6T Bx      ���'�   � � � �  nKH  <      ���'�   � � � �  @T =A      ���'�   � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �  LL F      ���k�  � � � �  |LL @@      ���k�  � � � �  LL  ?      ���k�  � � � �  |LL EE      ���+�  � � � �  LL AD      ���k�  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  }4T  x      ���  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �   x@5  x      ���  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �   LP* **      ��� ��  � � � �   I.. ..      ���  � � � �   M@& &&      �����  � � � �  H<& &&      �����  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �   MPI2 x      ��� ��  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  g2X2 x      ��� 	 � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �   _ M  x      ���+� 
 � � � �  _M  x      ���+�  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  2FI2 x      ��� ��  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  P M  x      ���	 
 � � � �  PM  x      ���	  � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �  @9  x      ���+�
  � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �  KH5  x      ���  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  }6T Bx      ���+�  � � � �  nKH  <      ���+�  � � � �  d@T =A      ���+�  � � � �  XDH =A      ���+�  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  _2X2 x      ����� 	 � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  _ M  x      ���+� 
 � � � �  _M  x      ���+�  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  }4T  x      ���  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  LL F      ���k�  � � � �  |LL @@      ���k�  � � � �  LL  ?      ���k�  � � � �  |LL EE      ���+�  � � � �  LL AD      ���k�  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �   ��	��
�B0                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    