pBAV       @� �� (  @  ������@   ����������@   ����������@   ����������@   ����������@   ����������@   ����������@   ����������@   ����������@   ����������@   ����������@   �������� ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  4        ���+�   � � � �  4        ���.�   � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �  d@V JJ      ����� 
 � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  7L F      ���k�  � � � �  |7L @@      ���k�  � � � �  7L  ?      ���k�  � � � �  |7L EE      ���+�  � � � �  7L AD      ���k�  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  lL> <      ���k�  � � � �  lL> 9;      ���k�  � � � �  lL>  8      ���k�  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  ,S MO      �����  � � � �  ,Y SV      �����  � � � �  ,] W      �����  � � � �  ,V PP      ���+�  � � � �  ,V QQ      ���+�  � � � �  ,V RR      ���+�  � � � �  ,S LL      ���  � � � �  ,S  K      �����  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  VS MO      �����  � � � �  VY SV      �����  � � � �  V] W      �����  � � � �  VV PP      ���+�  � � � �  VV QQ      ���+�  � � � �  VV RR      ���+�  � � � �  VS LL      ���  � � � �  VS  K      �����  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  2@R        ����� 	 � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  d O        ���  � � � �  }O        ���  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  2S  O      �����  � � � �  2Y SV      �����  � � � �  2] W      ���k�  � � � �  2V PR      ���+�  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  F@R        �����	 	 � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �  xPH        ���
  � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �  2S  O      �����_  � � � �  2Y SV      �����_  � � � �  2] W      �����_  � � � �  2V PR      �����_  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �   22V8���\D��X                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    