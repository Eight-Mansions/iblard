pBAV       �� ��   @  ������@�  ����������@�  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  N@V >>      �����   � � � �  U@_9@@      �����_   � � � �  P@^9AA      �����_   � � � �   U@[2CC      �����   � � � �   A@h;EE      �����   � � � �   @_ GG      �����   � � � �   @a HH      �����_   � � � �   S@k LL      �����   � � � �   Z@c MM      �����_   � � � �   n@f;JJ      �����  	 � � � �   P@q OO      �����   � � � �   <@w'QQ      �����   � � � �  #@o>SS      �����_   � � � �  7@r9TT      �����_   � � � �               �����_    � � � �               �����_    � � � �   Z@Z9<<      �����  � � � �   @n9>>      �����_  � � � �  d@^9@@      �����_ 
 � � � �   @_9AA      �����  � � � �   @f;CC      �����  � � � �  P@c9EE      �����_  � � � �   @e9GG      �����_  � � � �   4@X HH      �����  � � � �   4(Z JJ      �����  � � � �   4P\ LL      �����  � � � �  Z@k9MM      �����_  � � � �   Z@m9OO      �����  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �   F�Lj.��$z� �px\\�6Z��t	N�                                                                                                                                                                                                                                                                                                                                                                                                                                                                            