pBAV       �� ��   @  �����@   ���������@   ���������@   ���������@   ���������@   ���������@   ���������@   ���������@   ���������@   ���������@   ���������@   ���������@   ���������@   ���������@   ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    �������� \WF FF      ����KM   � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �  v2G  G      �����  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  i5T        ���k�  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  MT        ���  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  d@7        ���k�  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  f\H        ���+�  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  i O        �����  � � � �  iO        ���  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �   7@& &&      ����� 	 � � � �  2<& &&      ����� 	 � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  @9 99      ���+� 
 � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  U@E EE      ������	  � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �  FRH        ���+�
  � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �   U@7        �����  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  PPG  G      �����  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  n9T        �����  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �   n�p	P,  0�
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        