pBAV           ��   @  ����>@   ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  >    ��������  @<        �����   � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �   |                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            